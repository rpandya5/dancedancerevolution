// updated nov 18 10:46pm

module arrow_pattern_generator (
    input wire clock,                    // Clock input
    input wire reset,                    // Reset input
    input wire game_active,            // Signal from controller that game is in play state
    input wire beat_pulse,             // Timing pulse from audio/rhythm system
    
    // Arrow pattern outputs - active high when that arrow should be displayed
    output reg [3:0] pattern_out,      // Each bit represents an arrow (UDLR)
    output reg pattern_valid,          // High when pattern_out has valid data
    
    // Individual arrow creation signals
    output reg create_up,
    output reg create_down,
    output reg create_left,
    output reg create_right
);

    // Pattern definitions - 4'b(UDLR)
    localparam PATTERN_UP    = 4'b1000;
    localparam PATTERN_DOWN  = 4'b0100;
    localparam PATTERN_LEFT  = 4'b0010;
    localparam PATTERN_RIGHT = 4'b0001;
    
    // Valid pairs
    localparam PAIR_UP_DOWN   = 4'b1100;
    localparam PAIR_UP_LEFT   = 4'b1010;
    localparam PAIR_UP_RIGHT  = 4'b1001;
    localparam PAIR_DOWN_LEFT = 4'b0110;
    localparam PAIR_DOWN_RIGHT= 4'b0101;
    localparam PAIR_LEFT_RIGHT= 4'b0011;

    // LFSR for random pattern selection
    reg [15:0] lfsr;
    wire feedback = lfsr[15] ^ lfsr[14] ^ lfsr[12] ^ lfsr[3];

    // FSM states
    localparam IDLE     = 2'b00;
    localparam GENERATE = 2'b01;
    localparam HOLD    = 2'b10;
    
    reg [1:0] current_state;

    // Initialize with default values
    initial begin
        lfsr = 16'hACE1;  // Non-zero seed
        current_state = IDLE;
        pattern_valid = 0;
        pattern_out = 4'b0000;
        create_up = 0;
        create_down = 0;
        create_left = 0;
        create_right = 0;
    end

    // Combinational logic for setting create signals based on pattern_out
    always @(*) begin
        // Default all signals to 0
        create_up = 0;
        create_down = 0;
        create_left = 0;
        create_right = 0;

        if (pattern_valid) begin
            // Check each bit of pattern_out
            create_up = pattern_out[3];    // UDLR - bit 3 is up
            create_down = pattern_out[2];  // UDLR - bit 2 is down
            create_left = pattern_out[1];  // UDLR - bit 1 is left
            create_right = pattern_out[0]; // UDLR - bit 0 is right
        end
    end

    always @(posedge clock or posedge reset) begin
        if (reset) begin
            lfsr <= 16'hACE1;
            current_state <= IDLE;
            pattern_valid <= 0;
            pattern_out <= 4'b0000;
        end 
        else begin
            case (current_state)
                IDLE: begin
                    pattern_valid <= 0;
                    if (game_active && beat_pulse) begin
                        current_state <= GENERATE;
                    end
                end

                GENERATE: begin
                    // Update LFSR
                    lfsr <= {lfsr[14:0], feedback};
                    
                    // Use LFSR bits to determine pattern type and selection
                    case (lfsr[3:0])  // Use 4 bits for pattern selection
                        // Single arrows (4/16 chance = 25%)
                        4'b0000: pattern_out <= PATTERN_UP;
                        4'b0001: pattern_out <= PATTERN_DOWN;
                        4'b0010: pattern_out <= PATTERN_LEFT;
                        4'b0011: pattern_out <= PATTERN_RIGHT;
                        
                        // Pairs (12/16 chance = 75%)
                        4'b0100, 4'b0101: pattern_out <= PAIR_UP_DOWN;
                        4'b0110, 4'b0111: pattern_out <= PAIR_UP_LEFT;
                        4'b1000, 4'b1001: pattern_out <= PAIR_UP_RIGHT;
                        4'b1010, 4'b1011: pattern_out <= PAIR_DOWN_LEFT;
                        4'b1100, 4'b1101: pattern_out <= PAIR_DOWN_RIGHT;
                        4'b1110, 4'b1111: pattern_out <= PAIR_LEFT_RIGHT;
                    endcase
                    
                    pattern_valid <= 1;
                    current_state <= HOLD;
                end

                HOLD: begin
                    if (!beat_pulse) begin
                        current_state <= IDLE;
                        pattern_valid <= 0;
                    end
                end

                default: current_state <= IDLE;
            endcase
        end
    end
endmodule
